--------------------------------------------------------------------
-- Project     : DTP_Soundmachine
--
-- File Name   : Counter_Register.vhd
-- Description : 
--
--------------------------------------------------------------------
-- Change History

-- Date     |Name      |Modification
------------|----------|--------------------------------------------
-- 27.04.22 | rosraf   | creat file for pm2 project
--
--------------------------------------------------------------------